+incdir+${REPO_ROOT}/projects/myProjects${PROJECT_NUM}/src
./tb
