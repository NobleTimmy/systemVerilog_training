// Class: tb
//
// Top-level testbench, for the HELLO_WORLD project
module tb;
  initial begin
    $display("Hello World!");
    $finish;
  end
endmodule:tb
