+incdir+${REPO_ROOT}/projects/myProjects1/src
./tb